`ifndef STATE_SV
`define STATE_SV

int sequencer_finish = 0;
int driver_finish = 0;
int monitor_finish = 0;

`endif // STATE_SV
